module Datapath(
        input         clk, reset,
        input         memtoreg,
        input         dobranch,
        input         alusrcbimm,
        input  [4:0]  destreg,
        input         regwrite,
        input         jump,
        input  [2:0]  alucontrol,
        output        zero,
        output [31:0] pc,
        input  [31:0] instr,
        output [31:0] aluout,
        output [31:0] writedata,
        input  [31:0] readdata
);
        wire [31:0] pc, incpc;
        wire [31:0] signimm;
        wire [31:0] srca, srcb, srcbimm;
        wire [31:0] result;


        // Fetch: Reiche PC an Instruktionsspeicher weiter und update PC
        ProgramCounter pcenv(clk, reset, dobranch, signimm, jump, instr[25:0], pc, incpc);

        // Execute:
        // (a) Wähle Operanden aus
        SignExtension se(instr[15:0], signimm);
        assign srcbimm = alusrcbimm ? signimm : srcb;
        // (b) Führe Berechnung in der ALU durch
        ArithmeticLogicUnit alu((jump&&regwrite) ? incpc : srca,
                                 (jump&&regwrite) ? 32'b0 :srcbimm,
                                   alucontrol, aluout, zero);

        // (c) Wähle richtiges Ergebnis aus
        assign result = memtoreg ? readdata : aluout;

        // Memory: Datenwort das zur (möglichen) Speicherung an den Datenspeicher übertragen wird
        assign writedata = srcb;

        // Write-Back: Stelle Operanden bereit und schreibe das jeweilige Resultat zurück
        RegisterFile gpr(clk, regwrite, instr[25:21], instr[20:16],
                                   destreg, result, srca, srcb);

endmodule

module ProgramCounter(
        input         clk,
        input         reset,
        input         dobranch,
        input  [31:0] branchoffset,
        input         dojump,
        input  [25:0] jumptarget,
        output [31:0] progcounter,
        output [31:0] pc4
);
        reg  [31:0] pc;
        wire [31:0] incpc, branchpc, nextpc;

        // Inkrementiere Befehlszähler um 4 (word-aligned)
        Adder pcinc(.a(pc), .b(32'b100), .cin(1'b0), .y(incpc));
        // Berechne mögliches (PC-relatives) Sprungziel
        Adder pcbranch(.a(incpc), .b({branchoffset[29:0], 2'b00}), .cin(1'b0), .y(branchpc));
        // Wähle den nächsten Wert des Befehlszählers aus
        assign nextpc = dojump   ? {incpc[31:28], jumptarget, 2'b00} :
                                            dobranch ? branchpc :
                                                             incpc;
        // Der Befehlszähler ist ein Speicherbaustein
        always @(posedge clk)
        begin
                if (reset) begin // Initialisierung mit Adresse 0x00400000
                        pc <= 'h00400000;
                end else begin
                        pc <= nextpc;
                end
        end

        // Ausgabe
        assign progcounter = pc;
        assign pc4 = incpc;

endmodule

module RegisterFile(
	input         clk,
	input         we3,
	input  [4:0]  ra1, ra2, wa3,
	input  [31:0] wd3,
	output [31:0] rd1, rd2
);
	reg [31:0] registers[31:0];

	always @(posedge clk)
		if (we3) begin
			registers[wa3] <= wd3;
		end

	assign rd1 = (ra1 != 0) ? registers[ra1] : 0;
	assign rd2 = (ra2 != 0) ? registers[ra2] : 0;
endmodule

module Adder(
	input  [31:0] a, b,
	input         cin,
	output [31:0] y,
	output        cout
);
	assign {cout, y} = a + b + cin;
endmodule

module SignExtension(
	input  [15:0] a,
	output [31:0] y
);
	assign y = {{16{a[15]}}, a};
endmodule

module ArithmeticLogicUnit(
	input  [31:0] a, b,
	input  [2:0]  alucontrol,
	output [31:0] result,
	output        zero
);

reg [31:0] res;
reg z;

reg [63:0] mult;
wire [63:0] aext = {{32{1'b0}}, a};
wire [63:0] bext = {{32{1'b0}}, b};

always @(*)
    begin
        case(alucontrol)
            3'b000: res <= a < b ? 32'b1 : 32'b0;
            3'b001: res <= a - b;
            3'b101: res <= a + b;
            3'b110: res <= a | b;
            3'b111: res <= a & b;
            3'b010:
                begin
                    if (b != 32'b0)    // dann lui
                        res <= b << 16;
                    else
                        begin          //sonst ?
                            if (a == 32'b0)   // false bei bltz und 0 bei lui
                                res <= 32'b0;
                            else            // bltz a < 0
                                res <= a[31] == 1'b1 ? 32'b1 : 32'b0;

                        end
                end
            3'b100: mult <= aext * bext;
            3'b011: res <= b[1] == 1'b1 ? mult[31:0] : mult[63:32];
        endcase

        if(res == 32'b0)
            z = 1'b1;
        else
            z = 1'b0;
    end

assign result = res;
assign zero = z;

endmodule














